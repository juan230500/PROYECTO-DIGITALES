
// comparator2BitWithVHDL.v
module OR_GATE(
    input logic a, b,
    output logic c
);

assign c = a || b;
endmodule
